library ieee;
use ieee.std_logic_1164.all;

entity fetch is
    port(   clk         : in std_logic;
            instruction : in  std_logic_vector(0 to 31));

    
end entity fetch;